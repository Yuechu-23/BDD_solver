module test;
    rand bit [14:0] var_0;
    rand bit [12:0] var_1;
    rand bit [14:0] var_2;
    rand bit [7:0] var_3;
    rand bit [5:0] var_4;
    rand bit [11:0] var_5;
    rand bit [5:0] var_6;
    rand bit [11:0] var_7;
    rand bit [9:0] var_8;
    rand bit [10:0] var_9;
    rand bit [10:0] var_10;
    rand bit [10:0] var_11;
    rand bit [9:0] var_12;
    rand bit [3:0] var_13;
    rand bit [12:0] var_14;
    rand bit [14:0] var_15;
    rand bit [11:0] var_16;
    rand bit [12:0] var_17;
    rand bit [6:0] var_18;
    rand bit [6:0] var_19;
    rand bit [15:0] var_20;
    rand bit [3:0] var_21;
    rand bit [5:0] var_22;
    rand bit [13:0] var_23;
    rand bit [13:0] var_24;
    rand bit [12:0] var_25;
    rand bit [12:0] var_26;
    rand bit [8:0] var_27;
    rand bit [10:0] var_28;
    rand bit [12:0] var_29;
    rand bit [6:0] var_30;
    rand bit [7:0] var_31;
    rand bit [5:0] var_32;
    rand bit [13:0] var_33;
    rand bit [8:0] var_34;
    constraint cb {
        ~((~(var_13) * var_6));
        (var_10 != 16'h1a2);
        ((var_3 / 8'h5) - var_21);
        (var_31 | 8'h68);
        (~(var_22) | var_21);
        (var_11 ^ var_3);
        (!(~(var_24)) || var_32);
        (var_9 << 11'h4);
        ((var_32 + var_21) * 8'hf);
        (!(var_22) || var_1);
        (!(var_26) + 16'h1);
        (!(var_0) || var_19);
        (var_12 || var_14);
        (~(var_19) * var_6);
        (var_14 - 16'h160);
        (var_24 || var_10);
        ~((!(var_22) * var_13));
        (!(var_14) || var_23);
        ((var_31 != 8'h5d) * var_32);
        (!(var_2) | 1'h1);
        (var_20 << 16'hd);
        ((var_4 ^ var_22) - var_2);
        !(~((var_6 || var_17)));
        ((var_7 || var_17) || var_11);
        (!(var_16) != 16'h1);
        (var_13 - var_31);
        (var_31 || var_3);
        ((var_18 | 7'h2) * var_32);
        (var_6 >> 6'h3);
        ((var_3 * var_6) << 8'h2);
        (var_19 != var_7);
        (!(var_2) - 16'h0);
        (!(var_13) * var_31);
        ((!(var_33) || var_6) + var_34);
        !((~(var_1) >> 13'h2));
    }
endmodule
